-- Beau Bakken
-- University of Florida

library ieee;
use ieee.std_logic_1164.all;

package LC_3_PACKAGE is

constant WORD_SIZE : positive := 16;

end LC_3_PACKAGE;